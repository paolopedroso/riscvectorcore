    /*
     * Small Vector Floating Point RISC-V Core
     *
     * @copyright 2025 Paolo Pedroso <paoloapedroso@gmail.com>
     *
     * @license Apache 2.0
     *
     */

module top #(
    parameter int DATA_WIDTH = 32
) (
    input logic clk,
    input logic rst_n
);

// program_counter (
//     .clk(clk),
//     .rst_n(rst_n),
// );


endmodule
